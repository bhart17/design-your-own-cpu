module traffic_light_controller (
    output logic GREEN_LIGHT,
    output logic AMBER_LIGHT,
    output logic RED_LIGHT,
    input  logic BUTTON,
    input  logic clock,
    input  logic nreset
);

    timeunit 1ns; timeprecision 10ps;

    // Model your traffic light controller ASM here


endmodule
