module and2 (
    input  logic A,
    input  logic B,
    output logic Y
);

    timeunit 1ns; timeprecision 100ps;

    // Model the behaviour of the module here

    assign Y = A & B;

endmodule
